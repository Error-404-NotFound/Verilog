module four_level_nand_bench();
	reg a1;
	reg b1;
	reg c1;
	reg d1;
	wire y1;
	four_level_nand dUT_1(.a(a1),.b(b1),.c(c1),.d(d1),.y(y1));
	initial
	begin
		a1=1'b0;b1=1'b0;c1=1'b0;d1=1'b0;
	#100	a1=1'b0;b1=1'b0;c1=1'b0;d1=1'b1;
	#100	a1=1'b0;b1=1'b0;c1=1'b1;d1=1'b0;
	#100	a1=1'b0;b1=1'b0;c1=1'b1;d1=1'b1;
	#100	a1=1'b0;b1=1'b1;c1=1'b0;d1=1'b0;
	#100	a1=1'b0;b1=1'b1;c1=1'b0;d1=1'b1;
	#100	a1=1'b0;b1=1'b1;c1=1'b1;d1=1'b0;
	#100	a1=1'b0;b1=1'b1;c1=1'b1;d1=1'b1;
	#100	a1=1'b1;b1=1'b0;c1=1'b0;d1=1'b0;
	#100	a1=1'b1;b1=1'b0;c1=1'b0;d1=1'b1;
	#100	a1=1'b1;b1=1'b0;c1=1'b1;d1=1'b0;
	#100	a1=1'b1;b1=1'b0;c1=1'b1;d1=1'b1;
	#100	a1=1'b1;b1=1'b1;c1=1'b0;d1=1'b0;
	#100	a1=1'b1;b1=1'b1;c1=1'b0;d1=1'b1;
	#100	a1=1'b1;b1=1'b1;c1=1'b1;d1=1'b0;
	#100	a1=1'b1;b1=1'b1;c1=1'b1;d1=1'b1;
	end
endmodule