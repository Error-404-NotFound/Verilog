module OR(a,b,O);

	input a, b;
	output O; 
	assign O = a | b;

endmodule 